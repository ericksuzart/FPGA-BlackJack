// Made by: Erick

module Counter
#(parameter WIDTH = 12)
    (
        input clk_50M;              // 50 MHz clock
        input clk_2K;               // 2 kHz clock
        input i_Zero;               // Input para zerar o contador
        // -----------------------------------------------
        input i_Active;             // Input of 2sec from FSM
        input i_Reset;              // Input from reset push-button debouncer
        // -----------------------------------------------
        output [WIDTH-1:0] o_Count; // Saida do contador
        output o_TwoSec;            // Output indicates if 2 seconds elapsed
    );

    // Registrador para armazenar o numero do contador
    reg unsigned [WIDTH-1:0] r_Count;

    // Reset (i_Zero) if needed, or increment if i_Reset is enabled in high
    always @ (posedge clk_50M or posedge i_Zero)
    begin
        if (i_Zero)
            r_Count <= 0;
        else if (i_Reset == 1'b1)
            r_Count <= r_Count + 1;
    end

    // Increment if i_Active is enabled in high
    always @ (posedge clk_2k)
    begin
        if (i_Active == 1'b1 && r_Count < 2**(WIDTH) - 1)
            r_Count <= r_Count + 1;
        else if (r_Count == 2**(WIDTH) - 1)
            o_TwoSec <= 1;
    end

    assign o_Count = r_Count;
endmodule
